// hello.v : This file contains the 'top' module
module top;
 initial begin
    $display("Hello, world");
    $finish;
 end
endmodule

